module mod1(input a, b, c, d, s, output o);

    assign #10 w = ~a&~b&~c&~d | ~a&~b&~c&d | ~a&~b&c&~d | ~a&b&~c&d | ~a&b&c&~d |
        ~a&b&c&d | a&~b&~c&~d | a&~b&~c&d | a&~b&c&~d | a&b&c&~d ;

    assign #12 f = ~w&~b&c&~d | ~w&b&c&~d | w&~b&~c&~d | w&~b&~c&d |
        w&~b&c&~d | w&~b&c&d | w&b&c&~d | w&b&~c&d ;

    assign #14 g = ~a&~b&~c&~d | ~a&~b&c&d | ~a&b&~c&d | ~a&b&c&~d |
        ~a&b&c&d | a&~b&c&~d | a&~b&c&d | a&b&~c&d ;

    assign #5 o = s ? g : f;

endmodule